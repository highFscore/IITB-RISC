library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--library work;
--use MemoryComponent.all;



entity Memory is
  port(
    mem_out      : out std_logic_vector(15 downto 0);
    data         : in std_logic_vector(15 downto 0);
    addr         : in  std_logic_vector(15 downto 0);
    mem_write    : in  std_logic;
    clk          : in  std_logic
    );
end entity;


architecture Struct of Memory is
type MemArray is array(0 to 127) of std_logic_vector(15 downto 0);

constant INIT_MEMORY : MemArray := (
  0 => "0001000000010101",--adi(R0)
  1 => "0001001001010101",--adi(R1)
  2 => "1100000001010011",--lw(R2)
  3 => "0101010011010000",--sw
  4 => "0011011110101010",--lhi(R3)
  5 => "1001000001101010",--jlr()
  6 => "0000000000000000",
  7 => "0000000000000000",
  8 => "0000000000000000",
  9 => "0000000000000000",
  10 => "0000000000000000",
  11 => "0000000000000000",
  12 => "0000000000000000",
  13 => "0000000000000000",
  14 => "0000000000000000",
  15 => "1100001111000011",
  16 => "0000000000000000",
  17 => "0000000000000000",
  18 => "0000000000000000",
  19 => "0000000000000000",
  20 => "0000000000000000",
  21 => "0100101101001111",
  22 => "0000000000000000",
  23 => "0000000000000000",
  24 => "0000000000000000",
  25 => "0000000000000000",
  26 => "0000000000000000",
  27 => "0000000000000000",
  28 => "0000000000000000",
  29 => "0000000000000000",
  30 => "0000000000000000",
  31 => "0000000000000000",
  32 => "0000000000000000",
  33 => "0000000000000000",
  34 => "0000000000000000",
  35 => "0000000000000000",
  36 => "0000000000000000",
  37 => "0000000000000000",
  38 => "0000000000000000",
  39 => "0000000000000000",
  40 => "0000000000000000",
  41 => "0000000000000000",
  42 => "0000000000000000",
  43 => "0000000000000000",
  44 => "0000000000000000",
  45 => "0000000000000000",
  46 => "0000000000000000",
  47 => "0000000000000000",
  48 => "0000000000000000",
  49 => "0000000000000000",
  50 => "0000000000000000",
  51 => "0000000000000000",
  52 => "0000000000000000",
  53 => "0000000000000000",
  54 => "0000000000000000",
  55 => "0000000000000000",
  56 => "0000000000000000",
  57 => "0000000000000000",
  58 => "0000000000000000",
  59 => "0000000000000000",
  60 => "0000000000000000",
  61 => "0000000000000000",
  62 => "0000000000000000",
  63 => "0000000000000000",
  64 => "0000000000000000",
  65 => "0000000000000000",
  66 => "0000000000000000",
  67 => "0000000000000000",
  68 => "0000000000000000",
  69 => "0000000000000000",
  70 => "0000000000000000",
  71 => "0000000000000000",
  72 => "0000000000000000",
  73 => "0000000000000000",
  74 => "0000000000000000",
  75 => "0000000000000000",
  76 => "0000000000000000",
  77 => "0000000000000000",
  78 => "0000000000000000",
  79 => "0000000000000000",
  80 => "0000000000000000",
  81 => "0000000000000000",
  82 => "0000000000000000",
  83 => "0000000000000000",
  84 => "0000000000000000",
  85 => "0000000000000000",
  86 => "0000000000000000",
  87 => "0000000000000000",
  88 => "0000000000000000",
  89 => "0000000000000000",
  90 => "0000000000000000",
  91 => "0000000000000000",
  92 => "0000000000000000",
  93 => "0000000000000000",
  94 => "0000000000000000",
  95 => "0000000000000000",
  96 => "0000000000000000",
  97 => "0000000000000000",
  98 => "0000000000000000",
  99 => "0000000000000000",
  100 => "0000000000000000",
  101 => "0000000000000000",
  102 => "0000000000000000",
  103 => "0000000000000000",
  104 => "0000000000000000",
  105 => "0000000000000000",
  106 => "0000000000000000",
  107 => "0000000000000000",
  108 => "0000000000000000",
  109 => "0000000000000000",
  110 => "0000000000000000",
  111 => "0000000000000000",
  112 => "0000000000000000",
  113 => "0000000000000000",
  114 => "0000000000000000",
  115 => "0000000000000000",
  116 => "0000000000000000",
  117 => "0000000000000000",
  118 => "0000000000000000",
  119 => "0000000000000000",
  120 => "0000000000000000",
  121 => "0000000000000000",
  122 => "0000000000000000",
  123 => "0000000000000000",
  124 => "0000000000000000",
  125 => "0000000000000000",
  126 => "0000000000000000",
  127 => "0000000000000000"
);
  --signal memory_low : Memory;
  signal mem_array: MemArray := INIT_MEMORY;
  --signal addr_plus: std_logic_vector(15 downto 0);
begin
  --addr_plus <= std_logic_vector(unsigned(addr) + 1);
  process (clk) is
  begin
    if rising_edge(clk) then
      -- Write and bypass
      if mem_write = '1' then
        mem_array(to_integer(unsigned(addr(15 downto 0)))) <= data(15 downto 0);
        --mem_array(to_integer(unsigned(addr_plus(6 downto 0)))) <= data(15 downto 8);
      end if;

    end if;
  end process;

  mem_out(15 downto 0) <= mem_array(to_integer(unsigned(addr(6 downto 0))));
  --mem_out(7 downto 0) <= mem_array(to_integer(unsigned(addr(6 downto 0))));
end Struct;

